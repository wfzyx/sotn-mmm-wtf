pBAV        � �� f  @  ���� �8?   ���������8?   ���������8?   ���������8?   ���������8?   ���������8?   ���������8?   ���������8?   ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    ��������  �8    �������� A<         �����  � � � �  Z2<
        �����  � � � �  AH        �����  � � � �  Z2H
       �����  � � � �  AG        �����_  � � � �  Z2G
       �����_  � � � �  AG        �����  � � � �  Z2G
       �����  � � � �   @T        �����   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  x@T         �����_  � � � �  Z@T
        �����_  � � � �  x@T         �����_  � � � �  Z@T
        �����_  � � � �  x@T         �����_  � � � �  Z@T
        �����_  � � � �  x@T         �����_  � � � �  Z@T
        �����_  � � � �  x@T         �����_  � � � �  Z@T
        �����_  � � � �  x@T         �����_  � � � �  Z@T
        �����_  � � � �  x@T         �����_  � � � �  Z@T
        �����_  � � � �   x@T        �����  � � � �   Z@T
       �����  � � � �  x@YF x      �����_  � � � �  Z@YP x      �����_  � � � �               �����_  � � � �               �����_  � � � �  x@YF x      �����_  � � � �  Z@YP x      �����_  � � � �  x@T         �����_  � � � �  Z@T
        �����_  � � � �  x@T  x      �����_  � � � �  Z@T
 x      �����_  � � � �  x@T  x      �����_  � � � �  Z@T
 x      �����_  � � � �  x@YF x      �����_  � � � �  x@YP x      �����_  � � � �  x@T         �����_  � � � �  x@T
        �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T         �����_  � � � �  x@T
        �����_  � � � �  x@T         �����_  � � � �  x@T
        �����_  � � � �  x@T         �����_  � � � �  x@T
        �����_  � � � �  x@T         �����_  � � � �  x@T
        �����_  � � � �  x@T         �����_  � � � �  x@T
        �����_  � � � �  x@T         �����_  � � � �  x@T
        �����_  � � � �               �����_   � � � �               �����_   � � � �  x@T  x      �����_  � � � �  Z@T
 x      �����_  � � � �  x@T  x      �����_  � � � �  Z@T
 x      �����_  � � � �  x@YF x      �����_  � � � �  Z@YP x      �����_  � � � �  x@YF x      �����_  � � � �  Z@YP x      �����_  � � � �  x@T  x      �����_ 	 � � � �  Z@T
 x      �����_ 	 � � � �  x@T  x      �����_ 
 � � � �  Z@T
 x      �����_ 
 � � � �  x@T  x      �����_  � � � �  Z@T
 x      �����_  � � � �  x@T  x      �����  � � � �  Z@T  x      �����  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �               �����_  � � � �               �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �  x@TF       �����_  � � � �  x@TP       �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �  x@YF       �����  � � � �  Z@YP       �����  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �   R�x� �d�� �$v6nX�� ��b� �n                                                                                                                                                                                                                                                                                                                                                                                                                                                                               