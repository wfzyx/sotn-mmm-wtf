pBAV       0� �� `  @  ���� ��?�  �������� ��?�  ����������@�  ����������@�  ����������@�  ����������?�  ����������?�  ����������@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  @Rm       �����_  � � � �   @Rw       �����_  � � � �   @Rm       �����_  � � � �   @Rw       �����_  � � � �  @S;       �����  � � � �  @SE       �����_  � � � �   @R;       �����_  � � � �   @RE       �����_  � � � �  @S;       �����  � � � �  @SE       �����_  � � � �  @S;       �����  � � � �  @SE       �����_  � � � �  @S;       �����  � � � �  @SE       �����_  � � � �  @S;       �����  � � � �  @SE       �����_  � � � �  @S;       �����  � � � �  @SE       �����_  � � � �   @         �����_  � � � �   @         �����_  � � � �  @S;       ����� 	 � � � �  @SE       �����_ 	 � � � �  @S;       ����� 
 � � � �  @SE       �����_ 
 � � � �   @          �����_  � � � �   @          �����_  � � � �  @S;       �����  � � � �  @SE       �����_  � � � �  @S;       �����  � � � �  @SE       �����_  � � � �  @S;       �����  � � � �  @SE       �����_  � � � �  @S;       �����  � � � �  @SE       �����  � � � �   @Rm       �����  � � � �   @Rw       �����  � � � �  @S;       �����  � � � �  @SE       �����  � � � �  @S;       �����  � � � �  @SE       �����  � � � �    Q        �����_  � � � �    Q        �����_  � � � �    Q        �����_  � � � �    Q        �����_  � � � �    Q        �����_  � � � �    Q        �����_  � � � �  @NF       �����  � � � �  @NP       �����  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �   8������Fr�~�H�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                