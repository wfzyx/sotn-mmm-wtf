pBAV       �� ��	 �  @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �  x@T        �����_   � � � �  x@T
       �����_   � � � �  x@T        �����_   � � � �  Z@T
       �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �  x@MF       �����_   � � � �  Z@MP       �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        �����  � � � �  Z@T
       �����  � � � �  @H        ����� 
 � � � �  @H
       ����� 
 � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @Z9       �����  � � � �  @ZC       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@H        �����_  � � � �  Z@H
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@N9       �����_  � � � �  Z@NC       �����_  � � � �  x@Z9       �����_  � � � �  Z@ZC       �����_  � � � �  x@Z9       �����_  � � � �  Z@ZC       �����_  � � � �  x@Z9       �����  � � � �  Z@ZC       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@YF       �����_  � � � �  x@YP       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  @T  x      �����  � � � �  @T
 x      �����  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        ����� 	 � � � �  @T
       ����� 	 � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@T        �����  � � � �  Z@T
       �����_  � � � �  x@T        �����  � � � �  Z@T
       �����_  � � � �  x@T        ����� 	 � � � �  Z@T
       �����_ 	 � � � �     K        �����_  � � � �     K        �����_  � � � �  x@T        �����  � � � �  Z@T
       �����_  � � � �  x@T        �����  � � � �  Z@T
       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �   �v��\F�t�|h8� d�Hd.�`H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  