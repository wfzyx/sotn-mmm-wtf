pBAV       w �� J  @  ������?�  ����������?�  ����������?�  ����������?�  ��������
��?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �  @MF       �����   � � � �  Z@MP       �����   � � � �  @MF       �����  � � � �  Z@MP       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @H        �����  � � � �  Z@H
       �����  � � � �  @        �����  � � � �  @
       �����  � � � �  @$       �����  � � � �  @$
      �����  � � � �  @0 #      �����  � � � �  @0
#      �����  � � � �  @< $/      �����  � � � �  @<
$/      �����  � � � �  @H 0;      ����� 	 � � � �  @H
0;      ����� 	 � � � �  @T <G      �����  � � � �  @T
<G      �����  � � � �  @` HS      ����� 
 � � � �  @`
HS      ����� 
 � � � �  @l T_      �����  � � � �  n@l
T_      �����  � � � �  @        �����  � � � �  @
       �����  � � � �  @$       �����  � � � �  @$
      �����  � � � �  @0 #      �����  � � � �  @0
#      �����  � � � �  @< $/      �����  � � � �  @<
$/      �����  � � � �   @J 0;      �����  � � � �   @J
0;      �����  � � � �   @V <G      �����  � � � �   @V
<G      �����  � � � �   @b HS      �����  � � � �   @b
HS      �����  � � � �  @n T_      �����  � � � �  @n
T_      �����  � � � �   @K        �����  � � � �   @K
       �����  � � � �   @T        �����  � � � �   @T
       �����  � � � �  @AF       �����  � � � �  t@AP       �����  � � � �   @YF       �����  � � � �   @YP       �����  � � � �   @KF       �����  � � � �   @KP       �����  � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �               �����_   � � � �   �:(�j"�h�*�� H� �|�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            