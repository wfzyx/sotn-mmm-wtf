pBAV       �� �� 0  @  ������@�  ����������@�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �  @MF       �����   � � � �  Z@MP       �����   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        �����  � � � �  Z@T
       �����  � � � �  @H        �����  � � � �  Z@H
       �����  � � � �  @N9       �����  � � � �  @NC       �����  � � � �  @N9       �����  � � � �  @NC       �����  � � � �  @MF       �����  � � � �  Z@MP       �����  � � � �  @MF       �����  � � � �  Z@MP       �����  � � � �  @K        �����  � � � �  Z@K
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �   ���fvj�B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              