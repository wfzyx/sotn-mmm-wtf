pBAV       �� ��	 �  @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �   AK        �����  � � � �   2K
       �����  � � � �  AH        �����  � � � �  Z2H
       �����  � � � �  AG        �����_  � � � �  Z2G
       �����_  � � � �  AG        �����  � � � �  Z2G
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        �����  � � � �  @T
 x      �����  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @T        �����_  � � � �   @T
       �����_  � � � �   @T        �����_  � � � �   @T
       �����_  � � � �   @T        �����  � � � �   @T
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �  @P        �����  � � � �  n@P
       �����  � � � �   @K        �����  � � � �   @K        �����  � � � �  @P        �����_  � � � �  n@P
       �����_  � � � �  @P        �����  � � � �  n@P
       �����  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @Z        �����  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T  x      �����  � � � �  @T
 x      �����  � � � �  @T  x      �����  � � � �  @T
 x      �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        ����� 	 � � � �  @T
       ����� 	 � � � �   @T        �����  � � � �   @T
       �����  � � � �   @T        �����  � � � �   @T
       �����  � � � �   @T        �����  � � � �   @T
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        ����� 
 � � � �  @T
       ����� 
 � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �   R�x\� ^�z��`�D�`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            