pBAV       `� �� �  @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  �������� AH        �����   � � � �  Z2H
       �����   � � � �  AJ        �����   � � � �  Z2J
       �����   � � � �   AK        �����   � � � �   2K
       �����   � � � �  ZAMF       �����   � � � �  P2MP       �����   � � � �   AK        �����   � � � �   2K
       �����   � � � �   AK        �����   � � � �   2K
       �����   � � � �   AK        �����   � � � �   2K
       �����   � � � �   AK        �����   � � � �   2K
       �����   � � � �  AZ        �����  � � � �  Z2Z
       �����  � � � �  AU        �����  � � � �  Z2X
       �����  � � � �  AT        �����  � � � �  Z2T
       �����  � � � �  AY        �����  � � � �  Z2Y
       �����  � � � �  AS        �����  � � � �  Z2S
       �����  � � � �  AT        �����_  � � � �  Z2T
       �����_  � � � �  AT        �����_ 	 � � � �  Z2T
       �����_ 	 � � � �  AT        �����_ 
 � � � �  Z2T
       �����_ 
 � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@Y        �����_  � � � �  Z@Y
       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@Y        �����_  � � � �  Z@Y
       �����_  � � � �  x@Y        �����_  � � � �  Z@Y
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@YF        �����_  � � � �  Z@YP        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@YF x      �����_  � � � �  Z@YP x      �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@YF        �����_  � � � �  Z@YP        �����_  � � � �  x@YF        �����_  � � � �  Z@YP        �����_  � � � �  x@YF        �����_  � � � �  Z@YP        �����_  � � � �  x@M         �����  � � � �  Z@M
        �����  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   �� V�J@�>0�ZX��t&� �t�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                