pBAV       �� �� �  @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  �������� AH        �����   � � � �  Z2H
       �����   � � � �  AJ        �����   � � � �  Z2J
       �����   � � � �   AK        �����   � � � �   2K
       �����   � � � �  ZAMF       �����   � � � �  P2MP       �����   � � � �   AK        �����   � � � �   2K
       �����   � � � �   AK        �����   � � � �   2K
       �����   � � � �   AK        �����   � � � �   2K
       �����   � � � �   AK        �����   � � � �   2K
       �����   � � � �  AZ        �����  � � � �  Z2Z
       �����  � � � �  AU        �����  � � � �  Z2X
       �����  � � � �  AT        �����  � � � �  Z2T
       �����  � � � �  AY        �����  � � � �  Z2Y
       �����  � � � �  AS        �����  � � � �  Z2S
       �����  � � � �  AT        �����_  � � � �  Z2T
       �����_  � � � �  AT        �����_ 	 � � � �  Z2T
       �����_ 	 � � � �  AT        �����_ 
 � � � �  Z2T
       �����_ 
 � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����  � � � �  x@T
       �����  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  @Z        �����_  � � � �  n@Z
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  @Z        �����_  � � � �  n@Z
       �����_  � � � �  @Z        �����_  � � � �  n@Z
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@Z9       �����_  � � � �  Z@ZC       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@Z9       �����_  � � � �  Z@ZC       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@\9       �����_  � � � �  Z@\C       �����_  � � � �  x@X9       �����_  � � � �  Z@XC       �����_  � � � �  x@W9       �����_  � � � �  Z@WC       �����_  � � � �  x@M        �����  � � � �  Z@M
       �����  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   �� V�J@�>&� �t�&�� b�$�\                                                                                                                                                                                                                                                                                                                                                                                                                                                                              