pBAV       �� �� �  @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �   @K        �����  � � � �   @K
       �����  � � � �  @H        �����  � � � �  Z@H
       �����  � � � �  @G        �����_  � � � �  Z@G
       �����_  � � � �  @G        �����  � � � �  Z@G
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@Z9       �����_  � � � �  Z@ZC       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �    @K        �����_  � � � �    @K        �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �   @KF       �����_  � � � �   @KP       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K        �����_  � � � �  @T        �����_  � � � �  @T
       �����  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@T        �����_ 	 � � � �  Z@T
       �����_ 	 � � � �  x@T        �����_ 
 � � � �  Z@T
       �����_ 
 � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����  � � � �  Z@T        �����  � � � �  x@ZF       �����_  � � � �  Z@ZP       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@ZF       �����_  � � � �  Z@ZP       �����_  � � � �  x@TF       �����_  � � � �  x@TP       �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �  x@YF       �����_  � � � �  Z@YP       �����_  � � � �  x@YF       �����  � � � �  Z@YP       �����  � � � �   @T        �����  � � � �   @T
       �����  � � � �   @T        �����  � � � �   @T
       �����  � � � �   @T        �����_  � � � �   @T
       �����_  � � � �   @T        �����  � � � �   @T
       �����  � � � �   @T        �����_  � � � �   @T
       �����_  � � � �   @T        �����_  � � � �   @T
       �����_  � � � �   @T        �����_  � � � �   @T
       �����_  � � � �   @T        �����_  � � � �   @T
       �����_  � � � �   R�x� �d�� �$v6n� ��� �d.&�                                                                                                                                                                                                                                                                                                                                                                                                                                                                              