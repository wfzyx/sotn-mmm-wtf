pBAV       !  �� �  @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        �����  � � � �  Z@T
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             