pBAV       В �� l  @  ������?�  ����������?�  ����������@�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @Y        �����  � � � �  @Y
       �����  � � � �  @^C       �����  � � � �  Z@^M       �����  � � � �   @K         �����  � � � �   @K
        �����  � � � �  @T        �����  � � � �  @Tx       �����  � � � �  @T        �����  � � � �  @Tx       �����  � � � �  @T        �����  � � � �  @Tx       �����  � � � �              �����_   � � � �              �����_   � � � �              �����_   � � � �               �����_   � � � �  @T        �����  � � � �  @Tx       �����  � � � �  @T        �����  � � � �  @Tx       �����  � � � �  @T        ����� 	 � � � �  @Tx       ����� 	 � � � �  @T        ����� 
 � � � �  @Tx       ����� 
 � � � �  @T        �����  � � � �  @Tx       �����  � � � �  @T        �����  � � � �  @Tx       �����  � � � �  n@T        �����  � � � �  Z@T
       �����  � � � �   @K        �����_  � � � �   @K        �����_  � � � �   @KF       �����  � � � �   @KP       �����  � � � �   @KF       �����  � � � �   @KP       �����  � � � �   @KF       �����  � � � �   @KP       �����  � � � �   @KF       �����  � � � �   @KP       �����  � � � �   @YF       �����  � � � �   @YP       �����  � � � �   @YF       �����  � � � �   @YP       �����  � � � �   @YF       �����  � � � �   @YP       �����  � � � �   @KF       �����_  � � � �   @KP       �����_  � � � �  @T        �����_  � � � �  >Tx       �����_  � � � �   @T        �����_  � � � �   >T
       �����_  � � � �  @T        �����_  � � � �  >Tx       �����_  � � � �  @T        �����_  � � � �  >Tx       �����_  � � � �  @T        �����_  � � � �  >Tx       �����_  � � � �  @T        �����_ 
 � � � �  >Tx       �����_ 
 � � � �  @T        �����_  � � � �  >Tx       �����_  � � � �  @T        �����_  � � � �  >Tx       �����_  � � � �  @T        �����  � � � �  @Tx       �����  � � � �  @T        �����  � � � �  @Tx       �����  � � � �  @T        �����  � � � �  @Tx       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �   � \��n
~Z@
�
X&���>                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      