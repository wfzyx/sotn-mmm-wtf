pBAV       @�  �� P 
 @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  @T  x      �����  � � � �  Z@T
 x      �����  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_ 	 � � � �  Z@T
       �����_ 	 � � � �  x@R        �����_ 
 � � � �  Z@R
       �����_ 
 � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  @T        �����  � � � �  x@T
       �����  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   ��:�\dd� @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          