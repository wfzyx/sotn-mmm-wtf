pBAV       �B  �� �  @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        �����  � � � �  n@T
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        �����  � � � �  Z@T
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �   � ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        