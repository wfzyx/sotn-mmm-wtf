pBAV       @�  �� `  @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ����������@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@T        ����� 
 � � � �  P@T
       ����� 
 � � � �  x@T        �����  � � � �  Z@T
       �����  � � � �  x@O        �����  � � � �  Z@O
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����  � � � �  @T        �����  � � � �  @T        �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �   ��:�"PF\� �f�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    