pBAV        � ��	 �  @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @H        ����� 
 � � � �  Z@H
       ����� 
 � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@T        �����_  � � � �  x@T
       �����_  � � � �  x@T        �����_ 	 � � � �  x@T
       �����_ 	 � � � �  @YF       �����_  � � � �  n@YP       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@YF x      �����_  � � � �  Z@YP x      �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  @T        �����  � � � �  n@T
       �����  � � � �  @T        �����  � � � �  n@T
       �����  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  @T        �����_  � � � �  @T
       �����_  � � � �  @T        �����_  � � � �  @T
       �����_  � � � �  @T        �����_  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    T  x      �����  � � � �    T
 x      �����  � � � �    T  x      �����  � � � �    T
 x      �����  � � � �    T  x      �����  � � � �    T
 x      �����  � � � �    K        �����_  � � � �    K
       �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  @T        �����  � � � �  Z@T
       �����  � � � �  @T        �����  � � � �  Z@T
       �����  � � � �  @T        �����  � � � �  Z@T
       �����  � � � �   nbh6L��.�� ���"b`���<                                                                                                                                                                                                                                                                                                                                                                                                                                                                                