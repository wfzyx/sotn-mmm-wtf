pBAV       �� �� 2  @  ���� ��?�  �������� ��?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  @T        �����  � � � �   @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �   @T  x      �����  � � � �   @T
 x      �����_  � � � �  @T        ����� 
 � � � �  @T
       �����_ 
 � � � �  @T        ����� 	 � � � �  @T
       �����_ 	 � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @V        �����  � � � �  @V
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @T        �����  � � � �  @T
       �����_  � � � �  @V        �����  � � � �  @V
       �����_  � � � �   @<        �����  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �   @<        �����_  � � � �  x@ZF       �����  � � � �  Z@ZP       �����  � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �   H"�H:Z���l(��~�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        