pBAV       0� ��	 �  @  ������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ����������?�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  �������� @T        �����   � � � �  Z@T
       �����_   � � � �  @T        �����   � � � �  Z@T
       �����   � � � �  x@M        �����_  
 � � � �  Z@M
       �����_  
 � � � �  @T        �����   � � � �  Z@TP       �����_   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@T        �����_  � � � �  n@T
       �����_  � � � �  x@T        �����_  � � � �  n@T
       �����_  � � � �  x@O        �����  � � � �  n@O
       �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �     K        �����_  � � � �     K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �    K        �����_  � � � �    K
       �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �  @T        �����  � � � �  @T
       �����  � � � �   @K        �����_  � � � �   @K
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        ����� 	 � � � �  Z@T
       ����� 	 � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����  � � � �    K        �����  � � � �    K        �����  � � � �    K        �����  � � � �    K        �����  � � � �    K        �����  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �    K        �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  x@T        �����_  � � � �  Z@T
       �����_  � � � �  @T        �����  � � � �  Z@T
       �����  � � � �  @T        �����  � � � �  Z@T
       �����  � � � �  @T        �����  � � � �  Z@T
       �����  � � � �   j� fLbh6\��f��<��`�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    