pBAV        � ��    @  ������@�  ����������@�  ����������@�  ��������
��@�  ����������@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������   K        �����_    � � � �    K        �����_    � � � �    K        �����_    � � � �    K        �����_    � � � �    K        �����_    � � � �    K        �����_    � � � �    K        �����_    � � � �    K        �����_    � � � �  @MF       �����   � � � �  @MF
      �����   � � � �    K        �����_    � � � �    K        �����_    � � � �    K        �����_    � � � �    K        �����_    � � � �    K        �����_    � � � �    K        �����_    � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����   � � � �    K        �����   � � � �  @H        �����  � � � �  Z@H
       �����  � � � �   @S;       �����  � � � �   >SE       �����_  � � � �   @S;       �����  � � � �   >SE       �����_  � � � �  @N9       �����  � � � �  @NC       �����_  � � � �  @N9       �����  � � � �  @NC       �����_  � � � �  @N9       �����  � � � �  @NC       �����_  � � � �  @N9       ����� 	 � � � �  @NC       �����_ 	 � � � �  @S;       ����� 
 � � � �  @SE       �����_ 
 � � � �  @S;       �����  � � � �  @SE       �����_  � � � �   @N;       �����  � � � �   >NE       �����_  � � � �   @N;       �����  � � � �   >NE       �����_  � � � �  @N9       �����  � � � �  @NC       �����_  � � � �  @N9       �����  � � � �  @NC       �����_  � � � �   @N;       �����  � � � �   @NE       �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @H        �����  � � � �  x@H
       �����  � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �    K        �����_   � � � �   �|R �p�� �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        